module Traffic_Light ();
    
endmodule