module monitor_1001 (din, clk, rst_, find);
    input din, clk, rst_ ;
    output reg find;
    reg[3:0] shift_d4;
    reg[1:0] statur_timer;

    task satur;
        
    endtask
    
endmodule